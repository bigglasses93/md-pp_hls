//  /home/anh/workspace/mdg4a.r4257/src/bin/Linux-x86_64/gen_generic -n r2sqrt -f 0.5*sqrt(x) -b 26 -o 2 -w 7 -l 1.0 -r 2.0 -s 1 -z 1
//  sign : 1

module r2sqrt_0(input [6:0] adr, output reg [25:0] c);
  always_comb begin
    case (adr)
      7'h0: c = 26'h200ffc0;
      7'h1: c = 26'h202fdc3;
      7'h2: c = 26'h204f9cf;
      7'h3: c = 26'h206f3ea;
      7'h4: c = 26'h208ec19;
      7'h5: c = 26'h20ae262;
      7'h6: c = 26'h20cd6ca;
      7'h7: c = 26'h20ec957;
      7'h8: c = 26'h210ba0e;
      7'h9: c = 26'h212a8f4;
      7'ha: c = 26'h214960d;
      7'hb: c = 26'h2168161;
      7'hc: c = 26'h2186af2;
      7'hd: c = 26'h21a52c5;
      7'he: c = 26'h21c38e1;
      7'hf: c = 26'h21e1d48;
      7'h10: c = 26'h2200000;
      7'h11: c = 26'h221e10d;
      7'h12: c = 26'h223c074;
      7'h13: c = 26'h2259e38;
      7'h14: c = 26'h2277a5f;
      7'h15: c = 26'h22954ec;
      7'h16: c = 26'h22b2de3;
      7'h17: c = 26'h22d0549;
      7'h18: c = 26'h22edb21;
      7'h19: c = 26'h230af6f;
      7'h1a: c = 26'h2328238;
      7'h1b: c = 26'h234537e;
      7'h1c: c = 26'h2362346;
      7'h1d: c = 26'h237f194;
      7'h1e: c = 26'h239be6a;
      7'h1f: c = 26'h23b89cc;
      7'h20: c = 26'h23d53bf;
      7'h21: c = 26'h23f1c45;
      7'h22: c = 26'h240e361;
      7'h23: c = 26'h242a918;
      7'h24: c = 26'h2446d6c;
      7'h25: c = 26'h2463061;
      7'h26: c = 26'h247f1f9;
      7'h27: c = 26'h249b238;
      7'h28: c = 26'h24b7121;
      7'h29: c = 26'h24d2eb7;
      7'h2a: c = 26'h24eeafd;
      7'h2b: c = 26'h250a5f7;
      7'h2c: c = 26'h2525fa6;
      7'h2d: c = 26'h254180d;
      7'h2e: c = 26'h255cf31;
      7'h2f: c = 26'h2578512;
      7'h30: c = 26'h25939b5;
      7'h31: c = 26'h25aed1b;
      7'h32: c = 26'h25c9f48;
      7'h33: c = 26'h25e503e;
      7'h34: c = 26'h2600000;
      7'h35: c = 26'h261ae90;
      7'h36: c = 26'h2635bf1;
      7'h37: c = 26'h2650825;
      7'h38: c = 26'h266b32e;
      7'h39: c = 26'h2685d10;
      7'h3a: c = 26'h26a05cd;
      7'h3b: c = 26'h26bad66;
      7'h3c: c = 26'h26d53de;
      7'h3d: c = 26'h26ef938;
      7'h3e: c = 26'h2709d76;
      7'h3f: c = 26'h272409a;
      7'h40: c = 26'h273e2a6;
      7'h41: c = 26'h275839c;
      7'h42: c = 26'h277237f;
      7'h43: c = 26'h278c250;
      7'h44: c = 26'h27a6013;
      7'h45: c = 26'h27bfcc8;
      7'h46: c = 26'h27d9872;
      7'h47: c = 26'h27f3312;
      7'h48: c = 26'h280ccac;
      7'h49: c = 26'h2826541;
      7'h4a: c = 26'h283fcd2;
      7'h4b: c = 26'h2859362;
      7'h4c: c = 26'h28728f2;
      7'h4d: c = 26'h288bd85;
      7'h4e: c = 26'h28a511d;
      7'h4f: c = 26'h28be3ba;
      7'h50: c = 26'h28d7560;
      7'h51: c = 26'h28f060f;
      7'h52: c = 26'h29095c9;
      7'h53: c = 26'h2922491;
      7'h54: c = 26'h293b268;
      7'h55: c = 26'h2953f4f;
      7'h56: c = 26'h296cb49;
      7'h57: c = 26'h2985657;
      7'h58: c = 26'h299e07a;
      7'h59: c = 26'h29b69b5;
      7'h5a: c = 26'h29cf208;
      7'h5b: c = 26'h29e7976;
      7'h5c: c = 26'h2a00000;
      7'h5d: c = 26'h2a185a7;
      7'h5e: c = 26'h2a30a6e;
      7'h5f: c = 26'h2a48e55;
      7'h60: c = 26'h2a6115e;
      7'h61: c = 26'h2a7938b;
      7'h62: c = 26'h2a914dd;
      7'h63: c = 26'h2aa9555;
      7'h64: c = 26'h2ac14f5;
      7'h65: c = 26'h2ad93bf;
      7'h66: c = 26'h2af11b3;
      7'h67: c = 26'h2b08ed3;
      7'h68: c = 26'h2b20b21;
      7'h69: c = 26'h2b3869e;
      7'h6a: c = 26'h2b5014b;
      7'h6b: c = 26'h2b67b29;
      7'h6c: c = 26'h2b7f43b;
      7'h6d: c = 26'h2b96c80;
      7'h6e: c = 26'h2bae3fb;
      7'h6f: c = 26'h2bc5aad;
      7'h70: c = 26'h2bdd096;
      7'h71: c = 26'h2bf45b9;
      7'h72: c = 26'h2c0ba16;
      7'h73: c = 26'h2c22daf;
      7'h74: c = 26'h2c3a084;
      7'h75: c = 26'h2c51298;
      7'h76: c = 26'h2c683eb;
      7'h77: c = 26'h2c7f47e;
      7'h78: c = 26'h2c96453;
      7'h79: c = 26'h2cad36b;
      7'h7a: c = 26'h2cc41c7;
      7'h7b: c = 26'h2cdaf67;
      7'h7c: c = 26'h2cf1c4e;
      7'h7d: c = 26'h2d0887c;
      7'h7e: c = 26'h2d1f3f2;
      7'h7f: c = 26'h2d35eb1;
      default: c = 26'bx;
    endcase;
  end
endmodule // r2sqrt_0

//  /home/anh/workspace/mdg4a.r4257/src/bin/Linux-x86_64/gen_generic -n r2sqrt -f 0.5*sqrt(x) -b 26 -o 2 -w 7 -l 1.0 -r 2.0 -s 1 -z 1
//  sign : 1

module r2sqrt_1(input [6:0] adr, output reg [15:0] c);
  always_comb begin
    case (adr)
      7'h0: c = 16'hff80;
      7'h1: c = 16'hfe83;
      7'h2: c = 16'hfd89;
      7'h3: c = 16'hfc92;
      7'h4: c = 16'hfb9e;
      7'h5: c = 16'hfaac;
      7'h6: c = 16'hf9bd;
      7'h7: c = 16'hf8d1;
      7'h8: c = 16'hf7e7;
      7'h9: c = 16'hf700;
      7'ha: c = 16'hf61b;
      7'hb: c = 16'hf539;
      7'hc: c = 16'hf459;
      7'hd: c = 16'hf37b;
      7'he: c = 16'hf2a0;
      7'hf: c = 16'hf1c8;
      7'h10: c = 16'hf0f1;
      7'h11: c = 16'hf01d;
      7'h12: c = 16'hef4b;
      7'h13: c = 16'hee7b;
      7'h14: c = 16'hedad;
      7'h15: c = 16'hece1;
      7'h16: c = 16'hec17;
      7'h17: c = 16'heb4f;
      7'h18: c = 16'hea89;
      7'h19: c = 16'he9c5;
      7'h1a: c = 16'he903;
      7'h1b: c = 16'he843;
      7'h1c: c = 16'he785;
      7'h1d: c = 16'he6c9;
      7'h1e: c = 16'he60e;
      7'h1f: c = 16'he555;
      7'h20: c = 16'he49e;
      7'h21: c = 16'he3e8;
      7'h22: c = 16'he335;
      7'h23: c = 16'he282;
      7'h24: c = 16'he1d2;
      7'h25: c = 16'he123;
      7'h26: c = 16'he076;
      7'h27: c = 16'hdfca;
      7'h28: c = 16'hdf20;
      7'h29: c = 16'hde77;
      7'h2a: c = 16'hddd0;
      7'h2b: c = 16'hdd2a;
      7'h2c: c = 16'hdc85;
      7'h2d: c = 16'hdbe3;
      7'h2e: c = 16'hdb41;
      7'h2f: c = 16'hdaa1;
      7'h30: c = 16'hda02;
      7'h31: c = 16'hd965;
      7'h32: c = 16'hd8c9;
      7'h33: c = 16'hd82e;
      7'h34: c = 16'hd794;
      7'h35: c = 16'hd6fc;
      7'h36: c = 16'hd665;
      7'h37: c = 16'hd5cf;
      7'h38: c = 16'hd53b;
      7'h39: c = 16'hd4a7;
      7'h3a: c = 16'hd415;
      7'h3b: c = 16'hd384;
      7'h3c: c = 16'hd2f4;
      7'h3d: c = 16'hd266;
      7'h3e: c = 16'hd1d8;
      7'h3f: c = 16'hd14c;
      7'h40: c = 16'hd0c0;
      7'h41: c = 16'hd036;
      7'h42: c = 16'hcfad;
      7'h43: c = 16'hcf25;
      7'h44: c = 16'hce9e;
      7'h45: c = 16'hce18;
      7'h46: c = 16'hcd93;
      7'h47: c = 16'hcd0e;
      7'h48: c = 16'hcc8b;
      7'h49: c = 16'hcc09;
      7'h4a: c = 16'hcb88;
      7'h4b: c = 16'hcb08;
      7'h4c: c = 16'hca89;
      7'h4d: c = 16'hca0a;
      7'h4e: c = 16'hc98d;
      7'h4f: c = 16'hc911;
      7'h50: c = 16'hc895;
      7'h51: c = 16'hc81a;
      7'h52: c = 16'hc7a0;
      7'h53: c = 16'hc728;
      7'h54: c = 16'hc6af;
      7'h55: c = 16'hc638;
      7'h56: c = 16'hc5c2;
      7'h57: c = 16'hc54c;
      7'h58: c = 16'hc4d7;
      7'h59: c = 16'hc463;
      7'h5a: c = 16'hc3f0;
      7'h5b: c = 16'hc37e;
      7'h5c: c = 16'hc30c;
      7'h5d: c = 16'hc29b;
      7'h5e: c = 16'hc22b;
      7'h5f: c = 16'hc1bc;
      7'h60: c = 16'hc14d;
      7'h61: c = 16'hc0e0;
      7'h62: c = 16'hc072;
      7'h63: c = 16'hc006;
      7'h64: c = 16'hbf9a;
      7'h65: c = 16'hbf2f;
      7'h66: c = 16'hbec5;
      7'h67: c = 16'hbe5b;
      7'h68: c = 16'hbdf3;
      7'h69: c = 16'hbd8a;
      7'h6a: c = 16'hbd23;
      7'h6b: c = 16'hbcbc;
      7'h6c: c = 16'hbc56;
      7'h6d: c = 16'hbbf0;
      7'h6e: c = 16'hbb8b;
      7'h6f: c = 16'hbb27;
      7'h70: c = 16'hbac3;
      7'h71: c = 16'hba60;
      7'h72: c = 16'hb9fd;
      7'h73: c = 16'hb99c;
      7'h74: c = 16'hb93a;
      7'h75: c = 16'hb8da;
      7'h76: c = 16'hb87a;
      7'h77: c = 16'hb81a;
      7'h78: c = 16'hb7bb;
      7'h79: c = 16'hb75d;
      7'h7a: c = 16'hb6ff;
      7'h7b: c = 16'hb6a2;
      7'h7c: c = 16'hb645;
      7'h7d: c = 16'hb5e9;
      7'h7e: c = 16'hb58d;
      7'h7f: c = 16'hb532;
      default: c = 16'bx;
    endcase;
  end
endmodule // r2sqrt_1

//  /home/anh/workspace/mdg4a.r4257/src/bin/Linux-x86_64/gen_generic -n r2sqrt -f 0.5*sqrt(x) -b 26 -o 2 -w 7 -l 1.0 -r 2.0 -s 1 -z 1
//  sign : 1

module r2sqrt_2(input [6:0] adr, output reg [5:0] c);
  always_comb begin
    case (adr)
      7'h0: c = 6'h0;
      7'h1: c = 6'h1;
      7'h2: c = 6'h2;
      7'h3: c = 6'h3;
      7'h4: c = 6'h3;
      7'h5: c = 6'h4;
      7'h6: c = 6'h5;
      7'h7: c = 6'h5;
      7'h8: c = 6'h6;
      7'h9: c = 6'h7;
      7'ha: c = 6'h7;
      7'hb: c = 6'h8;
      7'hc: c = 6'h8;
      7'hd: c = 6'h9;
      7'he: c = 6'ha;
      7'hf: c = 6'ha;
      7'h10: c = 6'hb;
      7'h11: c = 6'hb;
      7'h12: c = 6'hc;
      7'h13: c = 6'hc;
      7'h14: c = 6'hd;
      7'h15: c = 6'hd;
      7'h16: c = 6'he;
      7'h17: c = 6'he;
      7'h18: c = 6'hf;
      7'h19: c = 6'hf;
      7'h1a: c = 6'h10;
      7'h1b: c = 6'h10;
      7'h1c: c = 6'h11;
      7'h1d: c = 6'h11;
      7'h1e: c = 6'h12;
      7'h1f: c = 6'h12;
      7'h20: c = 6'h12;
      7'h21: c = 6'h13;
      7'h22: c = 6'h13;
      7'h23: c = 6'h14;
      7'h24: c = 6'h14;
      7'h25: c = 6'h14;
      7'h26: c = 6'h15;
      7'h27: c = 6'h15;
      7'h28: c = 6'h16;
      7'h29: c = 6'h16;
      7'h2a: c = 6'h16;
      7'h2b: c = 6'h17;
      7'h2c: c = 6'h17;
      7'h2d: c = 6'h17;
      7'h2e: c = 6'h18;
      7'h2f: c = 6'h18;
      7'h30: c = 6'h18;
      7'h31: c = 6'h19;
      7'h32: c = 6'h19;
      7'h33: c = 6'h19;
      7'h34: c = 6'h1a;
      7'h35: c = 6'h1a;
      7'h36: c = 6'h1a;
      7'h37: c = 6'h1b;
      7'h38: c = 6'h1b;
      7'h39: c = 6'h1b;
      7'h3a: c = 6'h1c;
      7'h3b: c = 6'h1c;
      7'h3c: c = 6'h1c;
      7'h3d: c = 6'h1c;
      7'h3e: c = 6'h1d;
      7'h3f: c = 6'h1d;
      7'h40: c = 6'h1d;
      7'h41: c = 6'h1e;
      7'h42: c = 6'h1e;
      7'h43: c = 6'h1e;
      7'h44: c = 6'h1e;
      7'h45: c = 6'h1f;
      7'h46: c = 6'h1f;
      7'h47: c = 6'h1f;
      7'h48: c = 6'h1f;
      7'h49: c = 6'h20;
      7'h4a: c = 6'h20;
      7'h4b: c = 6'h20;
      7'h4c: c = 6'h20;
      7'h4d: c = 6'h21;
      7'h4e: c = 6'h21;
      7'h4f: c = 6'h21;
      7'h50: c = 6'h21;
      7'h51: c = 6'h21;
      7'h52: c = 6'h22;
      7'h53: c = 6'h22;
      7'h54: c = 6'h22;
      7'h55: c = 6'h22;
      7'h56: c = 6'h22;
      7'h57: c = 6'h23;
      7'h58: c = 6'h23;
      7'h59: c = 6'h23;
      7'h5a: c = 6'h23;
      7'h5b: c = 6'h24;
      7'h5c: c = 6'h24;
      7'h5d: c = 6'h24;
      7'h5e: c = 6'h24;
      7'h5f: c = 6'h24;
      7'h60: c = 6'h24;
      7'h61: c = 6'h25;
      7'h62: c = 6'h25;
      7'h63: c = 6'h25;
      7'h64: c = 6'h25;
      7'h65: c = 6'h25;
      7'h66: c = 6'h26;
      7'h67: c = 6'h26;
      7'h68: c = 6'h26;
      7'h69: c = 6'h26;
      7'h6a: c = 6'h26;
      7'h6b: c = 6'h26;
      7'h6c: c = 6'h27;
      7'h6d: c = 6'h27;
      7'h6e: c = 6'h27;
      7'h6f: c = 6'h27;
      7'h70: c = 6'h27;
      7'h71: c = 6'h27;
      7'h72: c = 6'h27;
      7'h73: c = 6'h28;
      7'h74: c = 6'h28;
      7'h75: c = 6'h28;
      7'h76: c = 6'h28;
      7'h77: c = 6'h28;
      7'h78: c = 6'h28;
      7'h79: c = 6'h28;
      7'h7a: c = 6'h29;
      7'h7b: c = 6'h29;
      7'h7c: c = 6'h29;
      7'h7d: c = 6'h29;
      7'h7e: c = 6'h29;
      7'h7f: c = 6'h29;
      default: c = 6'bx;
    endcase;
  end
endmodule // r2sqrt_2

